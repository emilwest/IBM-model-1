Ur v�gen  
 Sluta  
 Spring  Bis  
 Spring  
 Stanna h�r  
 Stoppa honom  
 Han kommer undan  
 Sl�pp mig  
 I konungens namn  
  Vad heter du  pojk  
  Dastan  sire  
 Och dina f�r�ldrar  
 Pojk  
  Bror  
 Ta med honom  
  R�rd av vad han s�g  
  adopterade kungen pojken  Dastan  till sin familj  
 En son utan kungligt blod  
 Och som inte tr�nade efter hans tron  
 Men det kanske var n�t annat som h�nde den dagen  
 N�t som var sv�rt att f�rst�  
 Dagen en pojke fr�n de mest ot�nkbaraste platserna   blev   en persisk prins  
15 �R SENARE 
 PERSISKA GR�NSOMR�DEN 
 DEN HELIGA STADEN ALAMUT 
  Mytiska Alamut  
 Vackrare �n jag trodde  
  Bli inte lurad  den �r som andra st�der  
 Veka l�nder ger veka m�n  
 De f�rr�dde oss och f�r nu betala  
 Vi f�r inte r�ra Alamut f�r far  
 Vissa betraktar den som helig  
 Men eftersom v�r vise far inte �r h�r s� ligger beslutet hos mig  
 En sista �verl�ggning med min nobla farbror och mina tv� br�der  
  Garsiv och  
 Var �r Dastan  
 Kom igen  
 Jag satsade hela min l�n  
 Det �r pinsamt  