st�ll konen p� den r�da kvadraten p� kvadraten
ta konen p� kvadraten
ta blocket
st�ll den r�da konen p� kvadraten
st�ll blocket p� den bl�a kvadraten p� kvadraten
st�ll den gr�na konen p� den bl�a cirkeln
st�ll den gr�na konen p� den r�da kvadraten
st�ll det bl�a blocket p� den r�da kvadraten
st�ll det r�da blocket p� den r�da kvadraten
st�ll den r�da konen p� den gr�na cirkeln p� kvadraten
ta den gr�na kuben p� den r�da cirkeln
ta den bl�a kuben p� den gr�na cirkeln
st�ll blocket p� cirkeln p� den r�da kvadraten
ta kuben
ta blocket
st�ll blocket p� cirkeln p� kvadraten
ta det gr�na blocket
ta kuben p� den r�da cirkeln
st�ll blocket p� den r�da kvadraten
st�ll blocket p� kvadraten p� den r�da cirkeln
ta kuben
st�ll den r�da konen p� kvadraten
st�ll kuben p� cirkeln p� den r�da cirkeln
st�ll det bl�a blocket p� den bl�a kvadraten
ta blocket p� kvadraten
ta det r�da blocket
ta den r�da kuben p� kvadraten
st�ll konen p� den r�da kvadraten p� den r�da kvadraten
st�ll blocket p� den r�da cirkeln
ta det gr�na blocket
st�ll blocket p� den r�da cirkeln
st�ll den bl�a kuben p� den r�da kvadraten
st�ll det bl�a blocket p� den bl�a kvadraten
ta konen
st�ll konen p� den r�da cirkeln p� kvadraten
ta det gr�na blocket
st�ll konen p� kvadraten p� den r�da kvadraten
st�ll kuben p� kvadraten p� cirkeln
ta blocket p� den r�da cirkeln
ta blocket
st�ll den r�da kuben p� den r�da kvadraten
ta det bl�a blocket
ta blocket
ta det gr�na blocket
st�ll den bl�a kuben p� kvadraten
st�ll blocket p� kvadraten p� den bl�a cirkeln
st�ll kuben p� den r�da cirkeln p� den r�da kvadraten
ta det r�da blocket
st�ll den bl�a kuben p� den gr�na cirkeln
st�ll det r�da blocket p� den bl�a cirkeln
st�ll kuben p� kvadraten
st�ll den bl�a konen p� kvadraten p� kvadraten
st�ll konen p� den r�da cirkeln p� kvadraten
st�ll det bl�a blocket p� den r�da cirkeln
st�ll kuben p� den r�da cirkeln p� cirkeln
ta kuben
st�ll den bl�a konen p� cirkeln
ta konen
st�ll den bl�a konen p� den r�da cirkeln p� kvadraten
st�ll den r�da kuben p� den r�da kvadraten
st�ll blocket p� den bl�a cirkeln
ta kuben p� cirkeln
st�ll kuben p� cirkeln p� cirkeln
st�ll blocket p� den r�da kvadraten
ta blocket p� cirkeln
st�ll det gr�na blocket p� den gr�na kvadraten
ta det r�da blocket
ta konen
st�ll kuben p� kvadraten
ta den r�da konen
st�ll konen p� kvadraten p� den r�da cirkeln
st�ll den r�da konen p� cirkeln
st�ll konen p� cirkeln p� den r�da cirkeln
ta det r�da blocket p� den bl�a kvadraten
ta det r�da blocket
ta blocket
st�ll det r�da blocket p� den gr�na cirkeln
st�ll blocket p� cirkeln p� cirkeln
st�ll konen p� cirkeln p� den r�da cirkeln
st�ll det r�da blocket p� cirkeln
st�ll konen p� kvadraten
st�ll blocket p� den bl�a kvadraten p� kvadraten
st�ll kuben p� den r�da cirkeln
ta det r�da blocket
st�ll det r�da blocket p� cirkeln p� den bl�a kvadraten
st�ll kuben p� den r�da kvadraten p� cirkeln
st�ll den bl�a konen p� den bl�a cirkeln
st�ll blocket p� kvadraten
st�ll kuben p� cirkeln
ta det gr�na blocket
st�ll den r�da konen p� kvadraten p� cirkeln
st�ll blocket p� den r�da cirkeln
st�ll den bl�a konen p� den r�da kvadraten
st�ll den r�da konen p� cirkeln
st�ll den bl�a konen p� den r�da cirkeln p� cirkeln
ta den bl�a konen
st�ll det r�da blocket p� den gr�na cirkeln
st�ll det gr�na blocket p� den r�da kvadraten
st�ll kuben p� den gr�na kvadraten
ta det bl�a blocket